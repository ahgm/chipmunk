module chipmunk

#include "/usr/include/chipmunk/chipmunk.h"
#flag -lchipmunk
